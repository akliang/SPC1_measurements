.option xbyname

* $HeadURL$
* $Id$

.subckt TAX
+ GLclamp
+ Vbias
+ VccSF
+ VccCSA
+ Vgnd
+ Val
+ Vreset
+ SFBgate
+ SFBgnd
+ SelGain
+ GlobRst1
+ GlobRst2
+ DLread1
+ DLread2
+ DLcap
+ DLgnd
+ DLrst1
+ DLrst2

.ends

.subckt G3
+ SAFT
+ SBEF
+ DGFLUSH
+ DGDATA
...
.ends

* Actual Setup:

xTAA TAX
+ PIN:
+ GLclamp=GLclamp
...

xG3C G3
+ SAFT=SAFT
+ SBEF=SBEF
+ DGDATA=DGDATA
...

* Voltages as generated by the PNC

VVout1  Vout1  0 0V
VVout2  Vout2  0 0V
VVout3  Vout3  0 0V
VVout4  Vout4  0 0V
VVout5  Vout5  0 0V
VVout6  Vout6  0 0V
VVout7  Vout7  0 0V
VVout8  Vout8  0 0V
VVout9  Vout9  0 0V
VVout10 Vout10 0 0V
VVout11 Vout11 0 0V
VVout12 Vout12 0 0V
VVout13 Vout13 0 0V
VVout14 Vout14 0 0V
VVout15 Vout15 0 0V
VVout16 Vout16 0 0V

* Primary functional mapping of Vout1..16

Vmap1x1  Vout1  Von      0V
Vmap2x1  Vout2  Voff     0V
Vmap3x1  Vout3  Qinj     0V
Vmap4x1  Vout4  Vref     0V
Vmap5x1  Vout5  VbiasNC  0V
Vmap6x1  Vout6  Vreset   0V
Vmap7x1  Vout7  VccCSA   0V
Vmap8x1  Vout8  VccSF    0V
Vmap9x1  Vout9  ValBgate PixLHI   0V
Vmap10x1 Vout10 VgndBgnd PixLLO   0V
Vmap11x1 Vout11 Spec1    DatLHI   0V
Vmap12x1 Vout12 Spec2    DatLLO   0V
Vmap13x1 Vout13 PixLLO   ValBgate 0V
Vmap14x1 Vout14 PixLHI   VgndBgnd 0V
Vmap15x1 Vout15 DatLLO   Spec1    0V
Vmap16x1 Vout16 DatLHI   Spec2    0V

* Additional mappings provided on PNC patchfield

Vmap2x2  Vout2  GLclamp  0V
Vmap4x2  Vout4  DLgndNC  0V
Vmap9x2  Vout9  Val       0V
Vmap9x3  Vout9  SFBgateNC 0V
Vmap10x2 Vout10 Vgnd      0V
Vmap10x3 Vout10 SFBgnd    0V
Vmap11x2 Vout11 VbiasNO   0V
Vmap11x3 Vout11 DLgndNO   0V
Vmap11x4 Vout11 DLcapNC   0V
Vmap12x2 Vout12 DLcapNO   0V
Vmap12x3 Vout12 SFBgateNO 0V
Vmap13x2 Vout13 SelgainNC 0V
Vmap13x3 Vout13 GlobRstNC 0V
Vmap14x2 Vout14 SelgainNO 0V
Vmap14x3 Vout14 GlobRstNO 0V
Vmap15x2 Vout15 DLreadNC  0V
Vmap15x3 Vout15 DLrstNC   0V
Vmap16x2 Vout16 DLreadNO  0V
Vmap16x3 Vout16 DLrstNO   0V

* Encode Current Limits in here, using some kind of spice syntax?

.subckt MAX333 SEL NC NO COMMON
Snc SEL NC COMMON NSW 17R 5pF
Sno SEL NO COMMON NSW 17R 5pF
.ends
VVVGND   GND 0 0V

Xu57ch3 G4IO5  Vout5  Vout11 Vbias      MAX333
* DLread1 shorted to DLread2 on the PNC
Xu57ch1 SAFT   Vout15 Vout16 DLread1    MAX333
* Xu57ch1 G4IO1  Vout15 Vout16 DLread1    MAX333
* Xu57ch2 DGDATA Vout13 Vout14 GlobRst    MAX333
Xu57ch2 G4IO2  Vout13 Vout14 GlobRst    MAX333
Xu57ch4	G4IO6  Vout13 Vout14 SelGain    MAX333

Xu56ch1 G4IO3  Vout15 Vout16 DLrst1     MAX333
Xu56ch2 G4IO4  Vout15 Vout16 DLrst2     MAX333
Xu56ch3 G4IO7  Vout11 Vout12 DLcap      MAX333
Xu56ch4 G4IO8  Vout9  Vout12 SFBgate    MAX333

* SMU mapping for TAA
Vsmu1x1  Vsmu1  Vout1    0V

Vsmu2x1  Vsmu2  Vout2    0V
Vsmu2x2  Vsmu2  Vout9    0V
Vsmu2x3  Vsmu2  Vout13   0V
* Vsmu2x4  Vsmu2  Vout15   0V
Vsmu2x5  Vsmu2  Vout5   0V
Vsmu2x6  Vsmu2  Vout7   0V
Vsmu2x7  Vsmu2  Vout10  0V
Vsmu2x8  Vsmu2  Vout11  0V
Vsmu2x9  Vsmu2  Vout12  0V

Vsmu3x1  Vsmu3  Vout3    0V

* Vsmu4x1  Vsmu4  Vout5    0V
* Vsmu4x3  Vsmu4  Vout13   0V
Vsmu4x4  Vsmu4  Vout15   0V

Vsmu5x1  Vsmu5  Vout6    0V
Vsmu5x2  Vsmu5  Vout4    0V

Vsmu6x1  Vsmu6  Vout8    0V

Vsmu7x1  Vsmu7  Vout14   0V

Vsmu8x1  Vsmu8  Vout16   0V

* SMU digio mapping
Vdigio1x1   CTRL10    0   0V
Vdigio1x2   CTRL9     0   0V
Vdigio1x3   PG5       0   0V
Vdigio1x4   PG4       0   0V
Vdigio1x5   PG3       0   0V
Vdigio1x6   SAFT      0   0V
Vdigio1x7   SBEF      0   0V
Vdigio1x8   IRST      0   0V
Vdigio1x9   PACLK     0   0V
Vdigio1x10  ABSEL     0   0V
Vdigio1x11  CTRL12    0   0V
Vdigio1x12  CTRL11    0   0V
Vdigio1x13  DG_EN     0   0V
Vdigio1x14  DG_CLK    0   0V
Vdigio2x1   DG_DATA   0   0V
Vdigio2x2   DG_FLSH   0   0V
Vdigio2x3   FAST_GATE 0   0V
Vdigio2x4   SYS_RSTb  0   0V

Vdigio2x5   G4IO10    0   0V
Vdigio2x6   G4IO9     0   0V
Vdigio2x7   G4IO6     0   0V
Vdigio2x8   G4IO5     0   0V
Vdigio2x9   G4IO2     0   0V

Vdigio2x10  G4IO3     0   0V
Vdigio2x11  G4IO4     0   0V
Vdigio2x12  G4IO7     0   0V
Vdigio2x13  G4IO8     0   0V
Vdigio2x14  G4IO1     0   0V





 
